library ieee;
use ieee.std_logic_1164.all;

package pwm_rom_pkg is
    constant PWM_LENGTH : integer := 2000;            -- rows in list
    subtype sample_t    is std_logic_vector(3 downto 0); -- Q4 Q3 Q2 Q1
    type rom_t          is array (0 to PWM_LENGTH-1) of sample_t;

    --  >>>  FULL PATTERN  (generated from your list)  <<<
    --  only six possible words appear: 0000, 0110, 0011, 0010, 0100, 1100
    constant PWM_ROM : rom_t := (
0    => "0000",
1    => "0110",
2    => "0110",
3    => "0110",
4    => "0110",
5    => "0110",
6    => "0110",
7    => "0110",
8    => "0110",
9    => "0110",
10   => "0110",
11   => "0110",
12   => "0011",
13   => "0110",
14   => "0110",
15   => "0110",
16   => "0110",
17   => "0110",
18   => "0110",
19   => "0110",
20   => "0110",
21   => "0110",
22   => "0110",
23   => "0010",
24   => "0011",
25   => "0010",
26   => "0110",
27   => "0110",
28   => "0110",
29   => "0110",
30   => "0110",
31   => "0110",
32   => "0110",
33   => "0110",
34   => "0110",
35   => "0011",
36   => "0011",
37   => "0011",
38   => "0110",
39   => "0110",
40   => "0110",
41   => "0110",
42   => "0110",
43   => "0110",
44   => "0110",
45   => "0110",
46   => "0010",
47   => "0011",
48   => "0011",
49   => "0011",
50   => "0010",
51   => "0110",
52   => "0110",
53   => "0110",
54   => "0110",
55   => "0110",
56   => "0110",
57   => "0110",
58   => "0010",
59   => "0011",
60   => "0011",
61   => "0011",
62   => "0010",
63   => "0110",
64   => "0110",
65   => "0110",
66   => "0110",
67   => "0110",
68   => "0110",
69   => "0110",
70   => "0011",
71   => "0011",
72   => "0011",
73   => "0011",
74   => "0011",
75   => "0110",
76   => "0110",
77   => "0110",
78   => "0110",
79   => "0110",
80   => "0110",
81   => "0010",
82   => "0011",
83   => "0011",
84   => "0011",
85   => "0011",
86   => "0011",
87   => "0010",
88   => "0110",
89   => "0110",
90   => "0110",
91   => "0110",
92   => "0110",
93   => "0011",
94   => "0011",
95   => "0011",
96   => "0011",
97   => "0011",
98   => "0011",
99   => "0011",
100  => "0110",
101  => "0110",
102  => "0110",
103  => "0110",
104  => "0010",
105  => "0011",
106  => "0011",
107  => "0011",
108  => "0011",
109  => "0011",
110  => "0011",
111  => "0011",
112  => "0010",
113  => "0110",
114  => "0110",
115  => "0110",
116  => "0010",
117  => "0011",
118  => "0011",
119  => "0011",
120  => "0011",
121  => "0011",
122  => "0011",
123  => "0011",
124  => "0010",
125  => "0110",
126  => "0110",
127  => "0110",
128  => "0011",
129  => "0011",
130  => "0011",
131  => "0011",
132  => "0011",
133  => "0011",
134  => "0011",
135  => "0011",
136  => "0011",
137  => "0110",
138  => "0110",
139  => "0110",
140  => "0011",
141  => "0011",
142  => "0011",
143  => "0011",
144  => "0011",
145  => "0011",
146  => "0011",
147  => "0011",
148  => "0011",
149  => "0010",
150  => "0110",
151  => "0010",
152  => "0011",
153  => "0011",
154  => "0011",
155  => "0011",
156  => "0011",
157  => "0011",
158  => "0011",
159  => "0011",
160  => "0011",
161  => "0010",
162  => "0110",
163  => "0010",
164  => "0011",
165  => "0011",
166  => "0011",
167  => "0011",
168  => "0011",
169  => "0011",
170  => "0011",
171  => "0011",
172  => "0011",
173  => "0010",
174  => "0110",
175  => "0011",
176  => "0011",
177  => "0011",
178  => "0011",
179  => "0011",
180  => "0011",
181  => "0011",
182  => "0011",
183  => "0011",
184  => "0011",
185  => "0011",
186  => "0110",
187  => "0011",
188  => "0011",
189  => "0011",
190  => "0011",
191  => "0011",
192  => "0011",
193  => "0011",
194  => "0011",
195  => "0011",
196  => "0011",
197  => "0011",
198  => "0010",
199  => "0011",
200  => "0011",
201  => "0011",
202  => "0011",
203  => "0011",
204  => "0011",
205  => "0011",
206  => "0011",
207  => "0011",
208  => "0011",
209  => "0011",
210  => "0010",
211  => "0011",
212  => "0011",
213  => "0011",
214  => "0011",
215  => "0011",
216  => "0011",
217  => "0011",
218  => "0011",
219  => "0011",
220  => "0011",
221  => "0011",
222  => "0010",
223  => "0011",
224  => "0011",
225  => "0011",
226  => "0011",
227  => "0011",
228  => "0011",
229  => "0011",
230  => "0011",
231  => "0011",
232  => "0011",
233  => "0011",
234  => "0010",
235  => "0011",
236  => "0011",
237  => "0011",
238  => "0011",
239  => "0011",
240  => "0011",
241  => "0011",
242  => "0011",
243  => "0011",
244  => "0011",
245  => "0011",
246  => "0010",
247  => "0011",
248  => "0011",
249  => "0011",
250  => "0011",
251  => "0011",
252  => "0011",
253  => "0011",
254  => "0011",
255  => "0011",
256  => "0011",
257  => "0011",
258  => "0010",
259  => "0011",
260  => "0011",
261  => "0011",
262  => "0011",
263  => "0011",
264  => "0011",
265  => "0011",
266  => "0011",
267  => "0011",
268  => "0011",
269  => "0011",
270  => "0010",
271  => "0011",
272  => "0011",
273  => "0011",
274  => "0011",
275  => "0011",
276  => "0011",
277  => "0011",
278  => "0011",
279  => "0011",
280  => "0011",
281  => "0011",
282  => "0010",
283  => "0011",
284  => "0011",
285  => "0011",
286  => "0011",
287  => "0011",
288  => "0011",
289  => "0011",
290  => "0011",
291  => "0011",
292  => "0011",
293  => "0011",
294  => "0010",
295  => "0011",
296  => "0011",
297  => "0011",
298  => "0011",
299  => "0011",
300  => "0011",
301  => "0011",
302  => "0011",
303  => "0011",
304  => "0011",
305  => "0011",
306  => "0010",
307  => "0011",
308  => "0011",
309  => "0011",
310  => "0011",
311  => "0011",
312  => "0011",
313  => "0011",
314  => "0011",
315  => "0011",
316  => "0011",
317  => "0011",
318  => "0110",
319  => "0011",
320  => "0011",
321  => "0011",
322  => "0011",
323  => "0011",
324  => "0011",
325  => "0011",
326  => "0011",
327  => "0011",
328  => "0011",
329  => "0010",
330  => "0110",
331  => "0011",
332  => "0011",
333  => "0011",
334  => "0011",
335  => "0011",
336  => "0011",
337  => "0011",
338  => "0011",
339  => "0011",
340  => "0011",
341  => "0010",
342  => "0110",
343  => "0010",
344  => "0011",
345  => "0011",
346  => "0011",
347  => "0011",
348  => "0011",
349  => "0011",
350  => "0011",
351  => "0011",
352  => "0011",
353  => "0110",
354  => "0110",
355  => "0010",
356  => "0011",
357  => "0011",
358  => "0011",
359  => "0011",
360  => "0011",
361  => "0011",
362  => "0011",
363  => "0011",
364  => "0011",
365  => "0110",
366  => "0110",
367  => "0110",
368  => "0011",
369  => "0011",
370  => "0011",
371  => "0011",
372  => "0011",
373  => "0011",
374  => "0011",
375  => "0011",
376  => "0010",
377  => "0110",
378  => "0110",
379  => "0110",
380  => "0010",
381  => "0011",
382  => "0011",
383  => "0011",
384  => "0011",
385  => "0011",
386  => "0011",
387  => "0011",
388  => "0110",
389  => "0110",
390  => "0110",
391  => "0110",
392  => "0010",
393  => "0011",
394  => "0011",
395  => "0011",
396  => "0011",
397  => "0011",
398  => "0011",
399  => "0011",
400  => "0110",
401  => "0110",
402  => "0110",
403  => "0110",
404  => "0110",
405  => "0011",
406  => "0011",
407  => "0011",
408  => "0011",
409  => "0011",
410  => "0011",
411  => "0010",
412  => "0110",
413  => "0110",
414  => "0110",
415  => "0110",
416  => "0110",
417  => "0010",
418  => "0011",
419  => "0011",
420  => "0011",
421  => "0011",
422  => "0011",
423  => "0110",
424  => "0110",
425  => "0110",
426  => "0110",
427  => "0110",
428  => "0110",
429  => "0010",
430  => "0011",
431  => "0011",
432  => "0011",
433  => "0011",
434  => "0010",
435  => "0110",
436  => "0110",
437  => "0110",
438  => "0110",
439  => "0110",
440  => "0110",
441  => "0110",
442  => "0011",
443  => "0011",
444  => "0011",
445  => "0011",
446  => "0010",
447  => "0110",
448  => "0110",
449  => "0110",
450  => "0110",
451  => "0110",
452  => "0110",
453  => "0110",
454  => "0010",
455  => "0011",
456  => "0011",
457  => "0011",
458  => "0110",
459  => "0110",
460  => "0110",
461  => "0110",
462  => "0110",
463  => "0110",
464  => "0110",
465  => "0110",
466  => "0110",
467  => "0011",
468  => "0011",
469  => "0010",
470  => "0110",
471  => "0110",
472  => "0110",
473  => "0110",
474  => "0110",
475  => "0110",
476  => "0110",
477  => "0110",
478  => "0110",
479  => "0010",
480  => "0011",
481  => "0110",
482  => "0110",
483  => "0110",
484  => "0110",
485  => "0110",
486  => "0110",
487  => "0110",
488  => "0110",
489  => "0110",
490  => "0110",
491  => "0110",
492  => "0010",
493  => "0110",
494  => "0110",
495  => "0110",
496  => "0110",
497  => "0110",
498  => "0110",
499  => "0110",
500  => "0110",
501  => "0110",
502  => "0110",
503  => "0110",
504  => "0100",
505  => "0110",
506  => "0110",
507  => "0110",
508  => "0110",
509  => "0110",
510  => "0110",
511  => "0110",
512  => "0110",
513  => "0110",
514  => "0110",
515  => "0100",
516  => "1100",
517  => "0110",
518  => "0110",
519  => "0110",
520  => "0110",
521  => "0110",
522  => "0110",
523  => "0110",
524  => "0110",
525  => "0110",
526  => "0110",
527  => "0100",
528  => "1100",
529  => "0100",
530  => "0110",
531  => "0110",
532  => "0110",
533  => "0110",
534  => "0110",
535  => "0110",
536  => "0110",
537  => "0110",
538  => "0110",
539  => "1100",
540  => "1100",
541  => "0100",
542  => "0110",
543  => "0110",
544  => "0110",
545  => "0110",
546  => "0110",
547  => "0110",
548  => "0110",
549  => "0110",
550  => "0100",
551  => "1100",
552  => "1100",
553  => "1100",
554  => "0100",
555  => "0110",
556  => "0110",
557  => "0110",
558  => "0110",
559  => "0110",
560  => "0110",
561  => "0110",
562  => "1100",
563  => "1100",
564  => "1100",
565  => "1100",
566  => "0100",
567  => "0110",
568  => "0110",
569  => "0110",
570  => "0110",
571  => "0110",
572  => "0110",
573  => "0100",
574  => "1100",
575  => "1100",
576  => "1100",
577  => "1100",
578  => "1100",
579  => "0110",
580  => "0110",
581  => "0110",
582  => "0110",
583  => "0110",
584  => "0110",
585  => "1100",
586  => "1100",
587  => "1100",
588  => "1100",
589  => "1100",
590  => "1100",
591  => "0100",
592  => "0110",
593  => "0110",
594  => "0110",
595  => "0110",
596  => "0100",
597  => "1100",
598  => "1100",
599  => "1100",
600  => "1100",
601  => "1100",
602  => "1100",
603  => "1100",
604  => "0110",
605  => "0110",
606  => "0110",
607  => "0110",
608  => "0100",
609  => "1100",
610  => "1100",
611  => "1100",
612  => "1100",
613  => "1100",
614  => "1100",
615  => "1100",
616  => "0110",
617  => "0110",
618  => "0110",
619  => "0110",
620  => "1100",
621  => "1100",
622  => "1100",
623  => "1100",
624  => "1100",
625  => "1100",
626  => "1100",
627  => "1100",
628  => "0100",
629  => "0110",
630  => "0110",
631  => "0100",
632  => "1100",
633  => "1100",
634  => "1100",
635  => "1100",
636  => "1100",
637  => "1100",
638  => "1100",
639  => "1100",
640  => "1100",
641  => "0110",
642  => "0110",
643  => "0100",
644  => "1100",
645  => "1100",
646  => "1100",
647  => "1100",
648  => "1100",
649  => "1100",
650  => "1100",
651  => "1100",
652  => "1100",
653  => "0110",
654  => "0110",
655  => "0100",
656  => "1100",
657  => "1100",
658  => "1100",
659  => "1100",
660  => "1100",
661  => "1100",
662  => "1100",
663  => "1100",
664  => "1100",
665  => "0100",
666  => "0110",
667  => "1100",
668  => "1100",
669  => "1100",
670  => "1100",
671  => "1100",
672  => "1100",
673  => "1100",
674  => "1100",
675  => "1100",
676  => "1100",
677  => "0100",
678  => "0100",
679  => "1100",
680  => "1100",
681  => "1100",
682  => "1100",
683  => "1100",
684  => "1100",
685  => "1100",
686  => "1100",
687  => "1100",
688  => "1100",
689  => "0100",
690  => "0100",
691  => "1100",
692  => "1100",
693  => "1100",
694  => "1100",
695  => "1100",
696  => "1100",
697  => "1100",
698  => "1100",
699  => "1100",
700  => "1100",
701  => "1100",
702  => "0100",
703  => "1100",
704  => "1100",
705  => "1100",
706  => "1100",
707  => "1100",
708  => "1100",
709  => "1100",
710  => "1100",
711  => "1100",
712  => "1100",
713  => "1100",
714  => "0100",
715  => "1100",
716  => "1100",
717  => "1100",
718  => "1100",
719  => "1100",
720  => "1100",
721  => "1100",
722  => "1100",
723  => "1100",
724  => "1100",
725  => "1100",
726  => "0100",
727  => "1100",
728  => "1100",
729  => "1100",
730  => "1100",
731  => "1100",
732  => "1100",
733  => "1100",
734  => "1100",
735  => "1100",
736  => "1100",
737  => "1100",
738  => "1100",
739  => "1100",
740  => "1100",
741  => "1100",
742  => "1100",
743  => "1100",
744  => "1100",
745  => "1100",
746  => "1100",
747  => "1100",
748  => "1100",
749  => "1100",
750  => "1100",
751  => "1100",
752  => "1100",
753  => "1100",
754  => "1100",
755  => "1100",
756  => "1100",
757  => "1100",
758  => "1100",
759  => "1100",
760  => "1100",
761  => "1100",
762  => "1100",
763  => "1100",
764  => "1100",
765  => "1100",
766  => "1100",
767  => "1100",
768  => "1100",
769  => "1100",
770  => "1100",
771  => "1100",
772  => "1100",
773  => "1100",
774  => "1100",
775  => "1100",
776  => "1100",
777  => "1100",
778  => "1100",
779  => "1100",
780  => "1100",
781  => "1100",
782  => "1100",
783  => "1100",
784  => "1100",
785  => "1100",
786  => "0100",
787  => "1100",
788  => "1100",
789  => "1100",
790  => "1100",
791  => "1100",
792  => "1100",
793  => "1100",
794  => "1100",
795  => "1100",
796  => "1100",
797  => "1100",
798  => "0100",
799  => "1100",
800  => "1100",
801  => "1100",
802  => "1100",
803  => "1100",
804  => "1100",
805  => "1100",
806  => "1100",
807  => "1100",
808  => "1100",
809  => "0100",
810  => "0100",
811  => "1100",
812  => "1100",
813  => "1100",
814  => "1100",
815  => "1100",
816  => "1100",
817  => "1100",
818  => "1100",
819  => "1100",
820  => "1100",
821  => "0100",
822  => "0100",
823  => "1100",
824  => "1100",
825  => "1100",
826  => "1100",
827  => "1100",
828  => "1100",
829  => "1100",
830  => "1100",
831  => "1100",
832  => "1100",
833  => "0100",
834  => "0110",
835  => "1100",
836  => "1100",
837  => "1100",
838  => "1100",
839  => "1100",
840  => "1100",
841  => "1100",
842  => "1100",
843  => "1100",
844  => "1100",
845  => "0110",
846  => "0110",
847  => "1100",
848  => "1100",
849  => "1100",
850  => "1100",
851  => "1100",
852  => "1100",
853  => "1100",
854  => "1100",
855  => "1100",
856  => "0100",
857  => "0110",
858  => "0110",
859  => "0100",
860  => "1100",
861  => "1100",
862  => "1100",
863  => "1100",
864  => "1100",
865  => "1100",
866  => "1100",
867  => "1100",
868  => "0100",
869  => "0110",
870  => "0110",
871  => "0100",
872  => "1100",
873  => "1100",
874  => "1100",
875  => "1100",
876  => "1100",
877  => "1100",
878  => "1100",
879  => "1100",
880  => "0110",
881  => "0110",
882  => "0110",
883  => "0110",
884  => "1100",
885  => "1100",
886  => "1100",
887  => "1100",
888  => "1100",
889  => "1100",
890  => "1100",
891  => "1100",
892  => "0110",
893  => "0110",
894  => "0110",
895  => "0110",
896  => "0100",
897  => "1100",
898  => "1100",
899  => "1100",
900  => "1100",
901  => "1100",
902  => "1100",
903  => "0100",
904  => "0110",
905  => "0110",
906  => "0110",
907  => "0110",
908  => "0100",
909  => "1100",
910  => "1100",
911  => "1100",
912  => "1100",
913  => "1100",
914  => "1100",
915  => "0110",
916  => "0110",
917  => "0110",
918  => "0110",
919  => "0110",
920  => "0110",
921  => "1100",
922  => "1100",
923  => "1100",
924  => "1100",
925  => "1100",
926  => "0100",
927  => "0110",
928  => "0110",
929  => "0110",
930  => "0110",
931  => "0110",
932  => "0110",
933  => "0100",
934  => "1100",
935  => "1100",
936  => "1100",
937  => "1100",
938  => "0100",
939  => "0110",
940  => "0110",
941  => "0110",
942  => "0110",
943  => "0110",
944  => "0110",
945  => "0110",
946  => "1100",
947  => "1100",
948  => "1100",
949  => "1100",
950  => "0110",
951  => "0110",
952  => "0110",
953  => "0110",
954  => "0110",
955  => "0110",
956  => "0110",
957  => "0110",
958  => "0100",
959  => "1100",
960  => "1100",
961  => "0100",
962  => "0110",
963  => "0110",
964  => "0110",
965  => "0110",
966  => "0110",
967  => "0110",
968  => "0110",
969  => "0110",
970  => "0110",
971  => "1100",
972  => "1100",
973  => "0110",
974  => "0110",
975  => "0110",
976  => "0110",
977  => "0110",
978  => "0110",
979  => "0110",
980  => "0110",
981  => "0110",
982  => "0110",
983  => "0100",
984  => "0100",
985  => "0110",
986  => "0110",
987  => "0110",
988  => "0110",
989  => "0110",
990  => "0110",
991  => "0110",
992  => "0110",
993  => "0110",
994  => "0110",
995  => "0110",
996  => "0110",
997  => "0110",
998  => "0110",
999  => "0110",
1000 => "0110",
1001 => "0110",
1002 => "0110",
1003 => "0110",
1004 => "0110",
1005 => "0110",
1006 => "0110",
1007 => "0010",
1008 => "0010",
1009 => "0110",
1010 => "0110",
1011 => "0110",
1012 => "0110",
1013 => "0110",
1014 => "0110",
1015 => "0110",
1016 => "0110",
1017 => "0110",
1018 => "0110",
1019 => "0010",
1020 => "0010",
1021 => "0110",
1022 => "0110",
1023 => "0110",
1024 => "0110",
1025 => "0110",
1026 => "0110",
1027 => "0110",
1028 => "0110",
1029 => "0110",
1030 => "0110",
1031 => "0011",
1032 => "0011",
1033 => "0010",
1034 => "0110",
1035 => "0110",
1036 => "0110",
1037 => "0110",
1038 => "0110",
1039 => "0110",
1040 => "0110",
1041 => "0110",
1042 => "0010",
1043 => "0011",
1044 => "0011",
1045 => "0010",
1046 => "0110",
1047 => "0110",
1048 => "0110",
1049 => "0110",
1050 => "0110",
1051 => "0110",
1052 => "0110",
1053 => "0110",
1054 => "0011",
1055 => "0011",
1056 => "0011",
1057 => "0011",
1058 => "0110",
1059 => "0110",
1060 => "0110",
1061 => "0110",
1062 => "0110",
1063 => "0110",
1064 => "0110",
1065 => "0010",
1066 => "0011",
1067 => "0011",
1068 => "0011",
1069 => "0011",
1070 => "0010",
1071 => "0110",
1072 => "0110",
1073 => "0110",
1074 => "0110",
1075 => "0110",
1076 => "0110",
1077 => "0011",
1078 => "0011",
1079 => "0011",
1080 => "0011",
1081 => "0011",
1082 => "0011",
1083 => "0110",
1084 => "0110",
1085 => "0110",
1086 => "0110",
1087 => "0110",
1088 => "0010",
1089 => "0011",
1090 => "0011",
1091 => "0011",
1092 => "0011",
1093 => "0011",
1094 => "0011",
1095 => "0010",
1096 => "0110",
1097 => "0110",
1098 => "0110",
1099 => "0110",
1100 => "0010",
1101 => "0011",
1102 => "0011",
1103 => "0011",
1104 => "0011",
1105 => "0011",
1106 => "0011",
1107 => "0010",
1108 => "0110",
1109 => "0110",
1110 => "0110",
1111 => "0110",
1112 => "0011",
1113 => "0011",
1114 => "0011",
1115 => "0011",
1116 => "0011",
1117 => "0011",
1118 => "0011",
1119 => "0011",
1120 => "0110",
1121 => "0110",
1122 => "0110",
1123 => "0010",
1124 => "0011",
1125 => "0011",
1126 => "0011",
1127 => "0011",
1128 => "0011",
1129 => "0011",
1130 => "0011",
1131 => "0011",
1132 => "0010",
1133 => "0110",
1134 => "0110",
1135 => "0010",
1136 => "0011",
1137 => "0011",
1138 => "0011",
1139 => "0011",
1140 => "0011",
1141 => "0011",
1142 => "0011",
1143 => "0011",
1144 => "0010",
1145 => "0110",
1146 => "0110",
1147 => "0011",
1148 => "0011",
1149 => "0011",
1150 => "0011",
1151 => "0011",
1152 => "0011",
1153 => "0011",
1154 => "0011",
1155 => "0011",
1156 => "0011",
1157 => "0110",
1158 => "0110",
1159 => "0011",
1160 => "0011",
1161 => "0011",
1162 => "0011",
1163 => "0011",
1164 => "0011",
1165 => "0011",
1166 => "0011",
1167 => "0011",
1168 => "0011",
1169 => "0110",
1170 => "0010",
1171 => "0011",
1172 => "0011",
1173 => "0011",
1174 => "0011",
1175 => "0011",
1176 => "0011",
1177 => "0011",
1178 => "0011",
1179 => "0011",
1180 => "0011",
1181 => "0010",
1182 => "0010",
1183 => "0011",
1184 => "0011",
1185 => "0011",
1186 => "0011",
1187 => "0011",
1188 => "0011",
1189 => "0011",
1190 => "0011",
1191 => "0011",
1192 => "0011",
1193 => "0010",
1194 => "0010",
1195 => "0011",
1196 => "0011",
1197 => "0011",
1198 => "0011",
1199 => "0011",
1200 => "0011",
1201 => "0011",
1202 => "0011",
1203 => "0011",
1204 => "0011",
1205 => "0010",
1206 => "0011",
1207 => "0011",
1208 => "0011",
1209 => "0011",
1210 => "0011",
1211 => "0011",
1212 => "0011",
1213 => "0011",
1214 => "0011",
1215 => "0011",
1216 => "0011",
1217 => "0010",
1218 => "0011",
1219 => "0011",
1220 => "0011",
1221 => "0011",
1222 => "0011",
1223 => "0011",
1224 => "0011",
1225 => "0011",
1226 => "0011",
1227 => "0011",
1228 => "0011",
1229 => "0011",
1230 => "0011",
1231 => "0011",
1232 => "0011",
1233 => "0011",
1234 => "0011",
1235 => "0011",
1236 => "0011",
1237 => "0011",
1238 => "0011",
1239 => "0011",
1240 => "0011",
1241 => "0011",
1242 => "0011",
1243 => "0011",
1244 => "0011",
1245 => "0011",
1246 => "0011",
1247 => "0011",
1248 => "0011",
1249 => "0011",
1250 => "0011",
1251 => "0011",
1252 => "0011",
1253 => "0011",
1254 => "0011",
1255 => "0011",
1256 => "0011",
1257 => "0011",
1258 => "0011",
1259 => "0011",
1260 => "0011",
1261 => "0011",
1262 => "0011",
1263 => "0011",
1264 => "0011",
1265 => "0011",
1266 => "0011",
1267 => "0011",
1268 => "0011",
1269 => "0011",
1270 => "0011",
1271 => "0011",
1272 => "0011",
1273 => "0011",
1274 => "0011",
1275 => "0011",
1276 => "0011",
1277 => "0010",
1278 => "0011",
1279 => "0011",
1280 => "0011",
1281 => "0011",
1282 => "0011",
1283 => "0011",
1284 => "0011",
1285 => "0011",
1286 => "0011",
1287 => "0011",
1288 => "0011",
1289 => "0010",
1290 => "0011",
1291 => "0011",
1292 => "0011",
1293 => "0011",
1294 => "0011",
1295 => "0011",
1296 => "0011",
1297 => "0011",
1298 => "0011",
1299 => "0011",
1300 => "0011",
1301 => "0010",
1302 => "0011",
1303 => "0011",
1304 => "0011",
1305 => "0011",
1306 => "0011",
1307 => "0011",
1308 => "0011",
1309 => "0011",
1310 => "0011",
1311 => "0011",
1312 => "0011",
1313 => "0010",
1314 => "0010",
1315 => "0011",
1316 => "0011",
1317 => "0011",
1318 => "0011",
1319 => "0011",
1320 => "0011",
1321 => "0011",
1322 => "0011",
1323 => "0011",
1324 => "0011",
1325 => "0110",
1326 => "0010",
1327 => "0011",
1328 => "0011",
1329 => "0011",
1330 => "0011",
1331 => "0011",
1332 => "0011",
1333 => "0011",
1334 => "0011",
1335 => "0011",
1336 => "0011",
1337 => "0110",
1338 => "0010",
1339 => "0011",
1340 => "0011",
1341 => "0011",
1342 => "0011",
1343 => "0011",
1344 => "0011",
1345 => "0011",
1346 => "0011",
1347 => "0011",
1348 => "0010",
1349 => "0110",
1350 => "0110",
1351 => "0011",
1352 => "0011",
1353 => "0011",
1354 => "0011",
1355 => "0011",
1356 => "0011",
1357 => "0011",
1358 => "0011",
1359 => "0011",
1360 => "0010",
1361 => "0110",
1362 => "0110",
1363 => "0010",
1364 => "0011",
1365 => "0011",
1366 => "0011",
1367 => "0011",
1368 => "0011",
1369 => "0011",
1370 => "0011",
1371 => "0011",
1372 => "0110",
1373 => "0110",
1374 => "0110",
1375 => "0010",
1376 => "0011",
1377 => "0011",
1378 => "0011",
1379 => "0011",
1380 => "0011",
1381 => "0011",
1382 => "0011",
1383 => "0011",
1384 => "0110",
1385 => "0110",
1386 => "0110",
1387 => "0110",
1388 => "0011",
1389 => "0011",
1390 => "0011",
1391 => "0011",
1392 => "0011",
1393 => "0011",
1394 => "0011",
1395 => "0010",
1396 => "0110",
1397 => "0110",
1398 => "0110",
1399 => "0110",
1400 => "0010",
1401 => "0011",
1402 => "0011",
1403 => "0011",
1404 => "0011",
1405 => "0011",
1406 => "0011",
1407 => "0110",
1408 => "0110",
1409 => "0110",
1410 => "0110",
1411 => "0110",
1412 => "0010",
1413 => "0011",
1414 => "0011",
1415 => "0011",
1416 => "0011",
1417 => "0011",
1418 => "0010",
1419 => "0110",
1420 => "0110",
1421 => "0110",
1422 => "0110",
1423 => "0110",
1424 => "0110",
1425 => "0011",
1426 => "0011",
1427 => "0011",
1428 => "0011",
1429 => "0011",
1430 => "0010",
1431 => "0110",
1432 => "0110",
1433 => "0110",
1434 => "0110",
1435 => "0110",
1436 => "0110",
1437 => "0010",
1438 => "0011",
1439 => "0011",
1440 => "0011",
1441 => "0011",
1442 => "0110",
1443 => "0110",
1444 => "0110",
1445 => "0110",
1446 => "0110",
1447 => "0110",
1448 => "0110",
1449 => "0110",
1450 => "0011",
1451 => "0011",
1452 => "0011",
1453 => "0010",
1454 => "0110",
1455 => "0110",
1456 => "0110",
1457 => "0110",
1458 => "0110",
1459 => "0110",
1460 => "0110",
1461 => "0110",
1462 => "0010",
1463 => "0011",
1464 => "0011",
1465 => "0110",
1466 => "0110",
1467 => "0110",
1468 => "0110",
1469 => "0110",
1470 => "0110",
1471 => "0110",
1472 => "0110",
1473 => "0110",
1474 => "0110",
1475 => "0011",
1476 => "0010",
1477 => "0110",
1478 => "0110",
1479 => "0110",
1480 => "0110",
1481 => "0110",
1482 => "0110",
1483 => "0110",
1484 => "0110",
1485 => "0110",
1486 => "0110",
1487 => "0010",
1488 => "0110",
1489 => "0110",
1490 => "0110",
1491 => "0110",
1492 => "0110",
1493 => "0110",
1494 => "0110",
1495 => "0110",
1496 => "0110",
1497 => "0110",
1498 => "0110",
1499 => "0000",
1500 => "0110",
1501 => "0110",
1502 => "0110",
1503 => "0110",
1504 => "0110",
1505 => "0110",
1506 => "0110",
1507 => "0110",
1508 => "0110",
1509 => "0110",
1510 => "0110",
1511 => "0100",
1512 => "0100",
1513 => "0110",
1514 => "0110",
1515 => "0110",
1516 => "0110",
1517 => "0110",
1518 => "0110",
1519 => "0110",
1520 => "0110",
1521 => "0110",
1522 => "0110",
1523 => "1100",
1524 => "0100",
1525 => "0110",
1526 => "0110",
1527 => "0110",
1528 => "0110",
1529 => "0110",
1530 => "0110",
1531 => "0110",
1532 => "0110",
1533 => "0110",
1534 => "0100",
1535 => "1100",
1536 => "1100",
1537 => "0110",
1538 => "0110",
1539 => "0110",
1540 => "0110",
1541 => "0110",
1542 => "0110",
1543 => "0110",
1544 => "0110",
1545 => "0110",
1546 => "1100",
1547 => "1100",
1548 => "1100",
1549 => "0100",
1550 => "0110",
1551 => "0110",
1552 => "0110",
1553 => "0110",
1554 => "0110",
1555 => "0110",
1556 => "0110",
1557 => "0100",
1558 => "1100",
1559 => "1100",
1560 => "1100",
1561 => "1100",
1562 => "0110",
1563 => "0110",
1564 => "0110",
1565 => "0110",
1566 => "0110",
1567 => "0110",
1568 => "0110",
1569 => "1100",
1570 => "1100",
1571 => "1100",
1572 => "1100",
1573 => "1100",
1574 => "0100",
1575 => "0110",
1576 => "0110",
1577 => "0110",
1578 => "0110",
1579 => "0110",
1580 => "0100",
1581 => "1100",
1582 => "1100",
1583 => "1100",
1584 => "1100",
1585 => "1100",
1586 => "1100",
1587 => "0110",
1588 => "0110",
1589 => "0110",
1590 => "0110",
1591 => "0110",
1592 => "0100",
1593 => "1100",
1594 => "1100",
1595 => "1100",
1596 => "1100",
1597 => "1100",
1598 => "1100",
1599 => "0100",
1600 => "0110",
1601 => "0110",
1602 => "0110",
1603 => "0110",
1604 => "1100",
1605 => "1100",
1606 => "1100",
1607 => "1100",
1608 => "1100",
1609 => "1100",
1610 => "1100",
1611 => "0100",
1612 => "0110",
1613 => "0110",
1614 => "0110",
1615 => "0100",
1616 => "1100",
1617 => "1100",
1618 => "1100",
1619 => "1100",
1620 => "1100",
1621 => "1100",
1622 => "1100",
1623 => "1100",
1624 => "0110",
1625 => "0110",
1626 => "0110",
1627 => "0100",
1628 => "1100",
1629 => "1100",
1630 => "1100",
1631 => "1100",
1632 => "1100",
1633 => "1100",
1634 => "1100",
1635 => "1100",
1636 => "0100",
1637 => "0110",
1638 => "0110",
1639 => "1100",
1640 => "1100",
1641 => "1100",
1642 => "1100",
1643 => "1100",
1644 => "1100",
1645 => "1100",
1646 => "1100",
1647 => "1100",
1648 => "0100",
1649 => "0110",
1650 => "0110",
1651 => "1100",
1652 => "1100",
1653 => "1100",
1654 => "1100",
1655 => "1100",
1656 => "1100",
1657 => "1100",
1658 => "1100",
1659 => "1100",
1660 => "0100",
1661 => "0110",
1662 => "0100",
1663 => "1100",
1664 => "1100",
1665 => "1100",
1666 => "1100",
1667 => "1100",
1668 => "1100",
1669 => "1100",
1670 => "1100",
1671 => "1100",
1672 => "1100",
1673 => "0110",
1674 => "0100",
1675 => "1100",
1676 => "1100",
1677 => "1100",
1678 => "1100",
1679 => "1100",
1680 => "1100",
1681 => "1100",
1682 => "1100",
1683 => "1100",
1684 => "1100",
1685 => "0110",
1686 => "1100",
1687 => "1100",
1688 => "1100",
1689 => "1100",
1690 => "1100",
1691 => "1100",
1692 => "1100",
1693 => "1100",
1694 => "1100",
1695 => "1100",
1696 => "1100",
1697 => "0100",
1698 => "1100",
1699 => "1100",
1700 => "1100",
1701 => "1100",
1702 => "1100",
1703 => "1100",
1704 => "1100",
1705 => "1100",
1706 => "1100",
1707 => "1100",
1708 => "1100",
1709 => "0100",
1710 => "1100",
1711 => "1100",
1712 => "1100",
1713 => "1100",
1714 => "1100",
1715 => "1100",
1716 => "1100",
1717 => "1100",
1718 => "1100",
1719 => "1100",
1720 => "1100",
1721 => "0100",
1722 => "1100",
1723 => "1100",
1724 => "1100",
1725 => "1100",
1726 => "1100",
1727 => "1100",
1728 => "1100",
1729 => "1100",
1730 => "1100",
1731 => "1100",
1732 => "1100",
1733 => "0100",
1734 => "1100",
1735 => "1100",
1736 => "1100",
1737 => "1100",
1738 => "1100",
1739 => "1100",
1740 => "1100",
1741 => "1100",
1742 => "1100",
1743 => "1100",
1744 => "1100",
1745 => "0100",
1746 => "1100",
1747 => "1100",
1748 => "1100",
1749 => "1100",
1750 => "1100",
1751 => "1100",
1752 => "1100",
1753 => "1100",
1754 => "1100",
1755 => "1100",
1756 => "1100",
1757 => "0100",
1758 => "1100",
1759 => "1100",
1760 => "1100",
1761 => "1100",
1762 => "1100",
1763 => "1100",
1764 => "1100",
1765 => "1100",
1766 => "1100",
1767 => "1100",
1768 => "1100",
1769 => "0100",
1770 => "1100",
1771 => "1100",
1772 => "1100",
1773 => "1100",
1774 => "1100",
1775 => "1100",
1776 => "1100",
1777 => "1100",
1778 => "1100",
1779 => "1100",
1780 => "1100",
1781 => "0100",
1782 => "1100",
1783 => "1100",
1784 => "1100",
1785 => "1100",
1786 => "1100",
1787 => "1100",
1788 => "1100",
1789 => "1100",
1790 => "1100",
1791 => "1100",
1792 => "1100",
1793 => "0100",
1794 => "1100",
1795 => "1100",
1796 => "1100",
1797 => "1100",
1798 => "1100",
1799 => "1100",
1800 => "1100",
1801 => "1100",
1802 => "1100",
1803 => "1100",
1804 => "1100",
1805 => "0100",
1806 => "1100",
1807 => "1100",
1808 => "1100",
1809 => "1100",
1810 => "1100",
1811 => "1100",
1812 => "1100",
1813 => "1100",
1814 => "1100",
1815 => "1100",
1816 => "1100",
1817 => "0110",
1818 => "1100",
1819 => "1100",
1820 => "1100",
1821 => "1100",
1822 => "1100",
1823 => "1100",
1824 => "1100",
1825 => "1100",
1826 => "1100",
1827 => "1100",
1828 => "1100",
1829 => "0110",
1830 => "0100",
1831 => "1100",
1832 => "1100",
1833 => "1100",
1834 => "1100",
1835 => "1100",
1836 => "1100",
1837 => "1100",
1838 => "1100",
1839 => "1100",
1840 => "0100",
1841 => "0110",
1842 => "0100",
1843 => "1100",
1844 => "1100",
1845 => "1100",
1846 => "1100",
1847 => "1100",
1848 => "1100",
1849 => "1100",
1850 => "1100",
1851 => "1100",
1852 => "0100",
1853 => "0110",
1854 => "0110",
1855 => "1100",
1856 => "1100",
1857 => "1100",
1858 => "1100",
1859 => "1100",
1860 => "1100",
1861 => "1100",
1862 => "1100",
1863 => "1100",
1864 => "0110",
1865 => "0110",
1866 => "0110",
1867 => "1100",
1868 => "1100",
1869 => "1100",
1870 => "1100",
1871 => "1100",
1872 => "1100",
1873 => "1100",
1874 => "1100",
1875 => "0100",
1876 => "0110",
1877 => "0110",
1878 => "0110",
1879 => "0100",
1880 => "1100",
1881 => "1100",
1882 => "1100",
1883 => "1100",
1884 => "1100",
1885 => "1100",
1886 => "1100",
1887 => "0100",
1888 => "0110",
1889 => "0110",
1890 => "0110",
1891 => "0100",
1892 => "1100",
1893 => "1100",
1894 => "1100",
1895 => "1100",
1896 => "1100",
1897 => "1100",
1898 => "1100",
1899 => "0110",
1900 => "0110",
1901 => "0110",
1902 => "0110",
1903 => "0110",
1904 => "1100",
1905 => "1100",
1906 => "1100",
1907 => "1100",
1908 => "1100",
1909 => "1100",
1910 => "0100",
1911 => "0110",
1912 => "0110",
1913 => "0110",
1914 => "0110",
1915 => "0110",
1916 => "0100",
1917 => "1100",
1918 => "1100",
1919 => "1100",
1920 => "1100",
1921 => "1100",
1922 => "0100",
1923 => "0110",
1924 => "0110",
1925 => "0110",
1926 => "0110",
1927 => "0110",
1928 => "0110",
1929 => "1100",
1930 => "1100",
1931 => "1100",
1932 => "1100",
1933 => "1100",
1934 => "0110",
1935 => "0110",
1936 => "0110",
1937 => "0110",
1938 => "0110",
1939 => "0110",
1940 => "0110",
1941 => "0100",
1942 => "1100",
1943 => "1100",
1944 => "1100",
1945 => "0100",
1946 => "0110",
1947 => "0110",
1948 => "0110",
1949 => "0110",
1950 => "0110",
1951 => "0110",
1952 => "0110",
1953 => "0110",
1954 => "1100",
1955 => "1100",
1956 => "1100",
1957 => "0110",
1958 => "0110",
1959 => "0110",
1960 => "0110",
1961 => "0110",
1962 => "0110",
1963 => "0110",
1964 => "0110",
1965 => "0110",
1966 => "0100",
1967 => "1100",
1968 => "0100",
1969 => "0110",
1970 => "0110",
1971 => "0110",
1972 => "0110",
1973 => "0110",
1974 => "0110",
1975 => "0110",
1976 => "0110",
1977 => "0110",
1978 => "0100",
1979 => "1100",
1980 => "0100",
1981 => "0110",
1982 => "0110",
1983 => "0110",
1984 => "0110",
1985 => "0110",
1986 => "0110",
1987 => "0110",
1988 => "0110",
1989 => "0110",
1990 => "0110",
1991 => "0100",
1992 => "0110",
1993 => "0110",
1994 => "0110",
1995 => "0110",
1996 => "0110",
1997 => "0110",
1998 => "0110",
1999 => "0110"
    );
end package;
